`timescale 1ns/1ps
/**********************************************************************************
 * net2axis verilog module                                                        *
 *                                                                                *
 * ISC License (ISC)                                                              *
 *                                                                                *
 * Copyright 2018 Lucas Brasilino <lucas.brasilino@gmail.com>                     *
 *                                                                                *
 * Refer to LICENSE file.                                                         *
 **********************************************************************************/

`ifndef DATAFILE
    `define DATAFILE ""
`endif

`define TO_STRING(s) `"s`"

module net2axis_tb;

    localparam C_TDATA_WIDTH = 32;

    localparam HALF_CORE_PERIOD = 5; // 100Mhz
    localparam PERIOD = HALF_CORE_PERIOD*2;
    localparam HARD_FINISH = 100;
    localparam INPUTFILE = `TO_STRING(`DATAFILE);
    localparam OUTPUTFILE = `TO_STRING(output.dat);
    reg                             ACLK;
    reg                             ARESETN;

    wire                            M_AXIS_TVALID;
    wire  [C_TDATA_WIDTH-1 : 0]     M_AXIS_TDATA;
    wire  [(C_TDATA_WIDTH/8)-1 : 0] M_AXIS_TKEEP;
    wire                            M_AXIS_TLAST;
    reg                             M_AXIS_TREADY;
    wire                            DONE;

    initial begin
        $timeformat(-9, 2, " ns", 20);
        ACLK = 1'b0;
        #(HALF_CORE_PERIOD);
        forever
            #(HALF_CORE_PERIOD) ACLK = ~ACLK;
    end

    initial begin
        ARESETN = 1'b0;
        #(PERIOD * 12);
        ARESETN = 1'b1;
    end

    initial begin
        wait (ARESETN == 1'b1);
        #(PERIOD * HARD_FINISH) $display("[%0t] Hard finish reached!",$time);
        $finish;
    end


    initial begin
        wait (DONE == 1'b1);
        #(PERIOD * 10);
        $display("[%0t] Simulation finished",$time);
        $finish;
    end

    wire clk;
    wire sync_rst;

    initial begin
        M_AXIS_TREADY = 1'b0;
        wait (sync_rst == 1'b1);
        #(PERIOD * 2);
        M_AXIS_TREADY = 1'b1;
    end

    net2axis_bd_wrapper DUT
        (.DONE(DONE),
            .M_AXIS_tdata(M_AXIS_TDATA),
            .M_AXIS_tkeep(M_AXIS_TKEEP),
            .M_AXIS_tlast(M_AXIS_TLAST),
            .M_AXIS_tready(M_AXIS_TREADY),
            .M_AXIS_tvalid(M_AXIS_TVALID),
            .clk(clk),
            .sync_rst(sync_rst));

    /*
    net2axis_master #(
        .C_INPUTFILE      (INPUTFILE),
        .C_TDATA_WIDTH    (C_TDATA_WIDTH   )
        ) net2axis (
        .ACLK             (ACLK            ),
        .ARESETN          (ARESETN         ),
        .DONE             (DONE            ),
        .M_AXIS_TVALID    (M_AXIS_TVALID   ),
        .M_AXIS_TDATA     (M_AXIS_TDATA    ),
        .M_AXIS_TKEEP     (M_AXIS_TKEEP    ),
        .M_AXIS_TLAST     (M_AXIS_TLAST    ),
        .M_AXIS_TREADY    (M_AXIS_TREADY));


    net2axis_slave #(
        .C_OUTPUTFILE   (OUTPUTFILE  ),
        .C_TDATA_WIDTH  (C_TDATA_WIDTH )
        ) net2axis_slave (
        .ACLK           (ACLK          ),
        .ARESETN        (ARESETN       ),
        .DONE           (DONE          ),
        .S_AXIS_TVALID  (M_AXIS_TVALID ),
        .S_AXIS_TDATA   (M_AXIS_TDATA  ),
        .S_AXIS_TKEEP   (M_AXIS_TKEEP  ),
        .S_AXIS_TLAST   (M_AXIS_TLAST  ),
        .S_AXIS_TREADY  (M_AXIS_TREADY ));
*/
endmodule
